module addressLatch(
input clk,
input[7:0] d,
input ce,
output reg[7:0] q
);
always @(posedge clk) begin
//just a big d flip flop 